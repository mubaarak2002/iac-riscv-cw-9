module CPU (


)(


);


endmodule